module ALU_Ctrl( funct_i, ALUOp_i, ALUCtrl_o );

//I/O ports
input      [6-1:0] funct_i;
input      [3-1:0] ALUOp_i;

output     [4-1:0] ALUCtrl_o;

//Internal Signals
reg        [4-1:0] ALUCtrl_o;

//Parameter

//Select exact operation

endmodule
